
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL; 
use IEEE.NUMERIC_STD.ALL;
use ieee.std_logic_unsigned.all;
use work.Fir_index_package.all;
use work.Package_FPDj.all;

entity Scope is
    generic(
        Horizontal_length : integer :=1280
    );
    port(
        Clk_i                               : in std_logic;
        Reset_i                             : in std_logic;      
        Audio_i                             : in std_logic_vector (15 downto 0); 
        Audio_Valid_i                       : in std_logic;  
        first_Row_i                         : in std_logic;     
        --BRAM Read interface
        clkb_i                              : IN STD_LOGIC;
        enb_i                               : IN STD_LOGIC;
        web_i                               : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
        addrb_i                             : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
        dinb_i                              : IN STD_LOGIC_VECTOR(30 DOWNTO 0);
        doutb_o                             : OUT STD_LOGIC_VECTOR(30 DOWNTO 0)
    );
end Scope;

architecture behevioral of Scope is

component blk_mem_gen_Scope IS
  PORT (
    clka    : IN STD_LOGIC;
    ena     : IN STD_LOGIC;
    wea     : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra   : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
    dina    : IN STD_LOGIC_VECTOR(30 DOWNTO 0);
    douta   : OUT STD_LOGIC_VECTOR(30 DOWNTO 0);
    clkb    : IN STD_LOGIC;
    enb     : IN STD_LOGIC;
    web     : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb   : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
    dinb    : IN STD_LOGIC_VECTOR(30 DOWNTO 0);
    doutb   : OUT STD_LOGIC_VECTOR(30 DOWNTO 0)
  );
END component;
      
signal Audio_amplitude_s    : std_logic_vector (30 downto 0);
signal Bram_write_EN        : std_logic_vector (0 downto 0);
signal Bram_Add_s           : std_logic_vector (10 DOWNTO 0);
signal din_s                : std_logic_vector (30 downto 0);
signal Audio_s              : std_logic_vector (15 downto 0); 
signal audio_downsample_counter : std_logic_vector (31 downto 0);
signal doutb_1s              : std_logic_vector (30 downto 0);
signal doutb_2s              : std_logic_vector (30 downto 0);
signal web_s                : std_logic_vector(0 downto 0);

begin       

-- convert audio from signed to unsigned
process ( Clk_i, Reset_i)
begin
    if Reset_i='1' then
        Audio_s <= (others=>'0');
    elsif rising_edge(Clk_i) then        
        Audio_s <=  not Audio_i(Audio_i'high) &  Audio_i(Audio_i'high- 1 downto 0);        
    end if;    
end process;
    
Audio_amplitude_s <="0000000000000000000000000000001" when Audio_s > (65535 -(2180*0)) else
                    "0000000000000000000000000000010" when Audio_s > (65535 -(2180*1)) else
                    "0000000000000000000000000000100" when Audio_s > (65535 -(2180*2)) else
                    "0000000000000000000000000001000" when Audio_s > (65535 -(2180*3)) else
                    "0000000000000000000000000010000" when Audio_s > (65535 -(2180*4)) else
                    "0000000000000000000000000100000" when Audio_s > (65535 -(2180*5)) else
                    "0000000000000000000000001000000" when Audio_s > (65535 -(2180*6)) else
                    "0000000000000000000000010000000" when Audio_s > (65535 -(2180*7)) else
                    "0000000000000000000000100000000" when Audio_s > (65535 -(2180*8)) else
                    "0000000000000000000001000000000" when Audio_s > (65535 -(2180*9)) else
                    "0000000000000000000010000000000" when Audio_s > (65535 -(2180*10)) else 
                    "0000000000000000000100000000000" when Audio_s > (65535 -(2180*11)) else 
                    "0000000000000000001000000000000" when Audio_s > (65535 -(2180*12)) else 
                    "0000000000000000010000000000000" when Audio_s > (65535 -(2180*13)) else 
                    "0000000000000000100000000000000" when Audio_s > (65535 -(2180*14)) else 
                    "0000000000000001000000000000000" when Audio_s > (65535 -(2180*15)) else 
                    "0000000000000010000000000000000" when Audio_s > (65535 -(2180*16)) else 
                    "0000000000000100000000000000000" when Audio_s > (65535 -(2180*17)) else 
                    "0000000000001000000000000000000" when Audio_s > (65535 -(2180*18)) else 
                    "0000000000010000000000000000000" when Audio_s > (65535 -(2180*19)) else 
                    "0000000000100000000000000000000" when Audio_s > (65535 -(2180*20)) else 
                    "0000000001000000000000000000000" when Audio_s > (65535 -(2180*21)) else 
                    "0000000010000000000000000000000" when Audio_s > (65535 -(2180*22)) else 
                    "0000000100000000000000000000000" when Audio_s > (65535 -(2180*23)) else                    
                    "0000001000000000000000000000000" when Audio_i > (65535 -(2180*24)) else                     
                    "0000010000000000000000000000000" when Audio_i > (65535 -(2180*25)) else 
                    "0000100000000000000000000000000" when Audio_i > (65535 -(2180*26)) else 
                    "0001000000000000000000000000000" when Audio_i > (65535 -(2180*27)) else 
                    "0010000000000000000000000000000" when Audio_i > (65535 -(2180*28)) else 
                    "0100000000000000000000000000000" when Audio_i > (65535 -(2180*29)) else 
                    "1000000000000000000000000000000" ;
                   





process ( Clk_i, Reset_i)
begin
    if Reset_i='1' then
    Bram_Add_s  <=(others=>'0');
     audio_downsample_counter <=(others=>'0');
    elsif rising_edge(Clk_i) then        
        if Audio_Valid_i = '1' then
           --audio_downsample_counter <= audio_downsample_counter+1;
            --if audio_downsample_counter= 37 then
            --    audio_downsample_counter <=(others=>'0');
                
                din_s <= Audio_amplitude_s;
                Bram_write_EN(0) <='1';
           
                if Bram_Add_s = Horizontal_length-1 then 
                    Bram_Add_s  <=(others=>'0');
                else
                    Bram_Add_s <= Bram_Add_s +1;
                end if;
            --end if;
        else
            Bram_write_EN(0) <='0'; 
        end if;
        
    end if;
end process;





--===================================
Blocl_Ram_Scope:blk_mem_gen_Scope
--===================================
  PORT map(
    clka    => Clk_i,                   
    ena     => '1',
    wea     => Bram_write_EN,         
    addra   => Bram_Add_s,            
    dina    => din_s,                 
    douta   => open,                  
    clkb    => clkb_i,   
    enb     => enb_i,    
    web     => "0",    
    addrb   => addrb_i,  
    dinb    => dinb_i,   
    doutb   => doutb_1s  
  );

  
--===================================
Blocl_Ram_Scope_saved :blk_mem_gen_Scope
--===================================
  PORT map(
    clka    => clkb_i,                   
    ena     => '0',
    wea     => "0",         
    addra   => Bram_Add_s,            
    dina    => din_s,                 
    douta   => open,                  
    clkb    => clkb_i,   
    enb     => enb_i,    
    web     => web_s,    
    addrb   => addrb_i,  
    dinb    => doutb_1s,   
    doutb   => doutb_2s  
  );
  doutb_o <= doutb_1s when first_Row_i='1' else doutb_2s;
  web_s <= "1" when first_Row_i='1' and web_i="1" else "0";

end behevioral;