-- Spec: 25 Hz to 20kHz
-- Sample frequency: 48kHz
-- Depth needed for min 4 samples at 20Hz: 2400*4= 9600

-- Depth to take 16384 or 8192

-- with FIR Depth at 16384 (2^14) and 16 bars:
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library work;
use work.Fir_index_package.all;



package Package_FPDj is


component Intensity_Bands_Extraction is
port(
    Clk_i                               : in std_logic;
    Reset_i                             : in std_logic;
    -- fft interface
    Frame_Index_i                       : in std_logic_vector (15 downto 0);
    Frame_start_i                       : in std_logic;
    Frame_end_i                         : in std_logic;
    Frame_Data_i                        : in std_logic_vector (31 downto 0);
    Frame_Data_valid_i                  : in std_logic;
    -- user Interface
    Bar_intensity_o                     : out  BarIndex_intensity_array;
    Data_Ready_o                        : out std_logic
);
end component;

component Intensity_Bands_Format is
port(
    Clk_i                               : in std_logic;
    Reset_i                             : in std_logic;      
    Bar_intensity_i                     : in  BarIndex_intensity_array;
    Data_Ready_i                        : in std_logic;
    Bar_intensity_o                     : out  BarIndex_intensity_array;
    Data_Ready_o                        : out std_logic    
);
end component;

 --------------------------------------------------------------------
 type Color_type is record    
        Red     : std_logic_vector(3 downto 0);
        Green   : std_logic_vector(3 downto 0);
        Blue    : std_logic_vector(3 downto 0);
end record;
    

 -- type BMP_array is array (0 to 163839) of std_logic_vector(11 downto 0);
-- constant FPDJ_Title :BMP_array:= (
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"777", x"ddd", x"fff", x"aaa", x"222",
    -- x"222", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"111", x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ddd", x"777", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"111", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"eee", x"888", x"111", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"555", x"aaa", x"ddd", x"ddd", x"ccc", x"555",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"333", x"bbb", x"fff", x"888", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"222",
    -- x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"222",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"888", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"555", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"555",
    -- x"ccc", x"fff", x"fff", x"fff", x"fff", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"111", x"ddd",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"aaa", x"333", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"666", x"aaa", x"888", x"555",
    -- x"777", x"bbb", x"eee", x"ddd", x"ccc", x"999", x"333", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"111", x"888", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"bbb", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"333", x"ccc", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"333", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"333", x"888", x"bbb", x"999", x"bbb", x"eee",
    -- x"ddd", x"888", x"bbb", x"eee", x"fff", x"fff", x"fff", x"eee",
    -- x"ccc", x"999", x"222", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"ccc", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"aaa", x"111", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa",
    -- x"333", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"444", x"aaa", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"eee", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"444", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"333",
    -- x"999", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"eee", x"444", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"999", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"eee", x"444", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ccc", x"eee", x"eee", x"888", x"111", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"777", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"999", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"222", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"444", x"bbb", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ccc", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"333", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"555", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"888",
    -- x"444", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"555",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"eee", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"eee", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"111", x"aaa", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"888", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"bbb", x"555", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"999", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"eee", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"111", x"999", x"eee", x"fff", x"eee",
    -- x"333", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"444", x"ddd", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"222", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc",
    -- x"222", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"444", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ccc", x"444", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"555", x"ddd", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"111", x"ddd", x"fff", x"fff", x"fff", x"fff",
    -- x"aaa", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"555", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"555", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"eee", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"888", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ddd", x"111", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"888", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"333",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"222", x"bbb", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"aaa", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"666", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"555", x"ccc", x"fff",
    -- x"777", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"333", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"ddd", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ccc", x"111", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"444", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"aaa", x"222", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"666", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"444", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"666", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"666", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"999", x"fff", x"fff", x"fff",
    -- x"eee", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"222",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"333", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"111",
    -- x"888", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ddd", x"222", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"555", x"eee", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"888", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"888",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"bbb", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"333", x"ddd", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"444", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"ccc",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"999",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999",
    -- x"000", x"000", x"777", x"ddd", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"333", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"888",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"555", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"222", x"ccc",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"555", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"666", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"bbb", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"444", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"777", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"aaa", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"555", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"777", x"000", x"000", x"000", x"666", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ddd", x"111", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"888", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"222", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"444", x"eee", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ccc", x"222", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"aaa", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"555", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"777", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"777", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"eee", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"111", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"555", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"555", x"000", x"000", x"000", x"555", x"eee", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"888", x"ddd", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"777",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"888", x"ddd", x"fff",
    -- x"fff", x"ccc", x"222", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"bbb", x"111", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"777",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"888", x"000", x"000", x"000", x"000", x"000", x"000", x"222",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"333",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"888", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"222", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"aaa", x"888", x"666", x"666",
    -- x"888", x"888", x"222", x"000", x"555", x"bbb", x"fff", x"fff",
    -- x"fff", x"fff", x"ccc", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"222", x"000", x"000", x"000", x"444", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"111", x"444", x"777",
    -- x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"222", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"555", x"eee", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"888", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"666", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"888",
    -- x"000", x"888", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"666", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"ddd",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"444", x"000", x"000", x"000", x"000", x"000", x"000", x"555",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"111", x"ddd",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"888", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"666", x"111", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"222", x"999",
    -- x"eee", x"fff", x"555", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"444", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ccc", x"000", x"000", x"000", x"000", x"333",
    -- x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"666",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"666", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"999", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"555", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"777", x"000",
    -- x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ddd", x"333", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"777", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"111",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"bbb", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"666", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"666",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"222", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"777", x"000", x"000", x"000", x"000",
    -- x"111", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee",
    -- x"333", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"999",
    -- x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"222", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"888", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"444", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"555", x"111", x"ccc",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"ddd", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"888", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"666", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"444", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"ddd", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"333", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"eee", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ddd", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"888", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"333",
    -- x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"444", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"222", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"555", x"000", x"bbb", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"555", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"777", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"555",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"111", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"222", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"666", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"444", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"777", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"999", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"777", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"111",
    -- x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"111", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"333", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"555", x"000", x"333", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"aaa", x"111", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ddd", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"666",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ccc", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"999", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"444", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"666", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"777", x"000",
    -- x"000", x"222", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"111",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"111", x"ddd", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"aaa", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"777",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"777", x"000", x"000", x"333", x"fff", x"fff",
    -- x"fff", x"fff", x"ccc", x"444", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"888",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ccc", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"444", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"eee", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"111", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"444", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"222", x"000",
    -- x"000", x"000", x"000", x"333", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"333", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"999", x"000", x"000", x"000", x"000", x"999", x"ccc",
    -- x"aaa", x"555", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"ddd", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"999",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"eee", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"ddd", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"444", x"bbb", x"eee", x"fff", x"fff",
    -- x"ddd", x"444", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"666", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"222", x"eee", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"666", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"ddd", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"444", x"ccc", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"aaa", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"333", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"666", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ddd", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"aaa",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"111", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"bbb", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"333", x"eee", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ccc", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"666", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"111", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"555", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"444", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"222", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"666",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"666", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"999", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"666", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"ccc", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"444", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"ddd", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"222", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"ccc",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"555", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"555", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"999", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"111", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ccc", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"111", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"555", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"888",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"444", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"666", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"111", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"222", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"777", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"555", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"ddd",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"222", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"666", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"555", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"999", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ccc", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"888", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ccc", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"222", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"777", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"bbb", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"999", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"888",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ddd", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"777",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"555", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"ccc",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"333", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"aaa",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"666", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"888", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"777", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"eee", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"444", x"eee", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"444", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"444", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"555",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"333", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"111", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"aaa",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"aaa",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"bbb", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"111", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"444", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"555", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"444", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"333", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"111", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"333", x"ddd", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"111", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"eee", x"666", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"888", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"555",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"bbb",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"555", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"777", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"999", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"666", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"eee", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"555", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"222", x"ddd", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"222", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"555", x"ccc", x"eee",
    -- x"fff", x"fff", x"eee", x"999", x"111", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"777",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"444", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"ddd",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"555", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"444", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"888", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"333", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"333",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"bbb", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"999", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"777", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"333", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"222", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"555", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"222", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"111", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"222", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"777",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"333", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"111", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"666",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"777", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"777", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"888", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"eee", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"333",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ccc", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"ddd", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"555", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"333",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"111", x"ddd", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ccc", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"222",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"222", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"777", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"777", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"999",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"111", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"111", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ccc", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"555", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"111", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"ddd", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"666", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"888", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"888", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"555", x"000", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"666",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"222", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"bbb",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ccc", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"555", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"333",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"111", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"bbb", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"555", x"000", x"222", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"444", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"999", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"555", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"555", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"999",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"ddd", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"666", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"888", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"888", x"000", x"000", x"777", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"777", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"111", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"111", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"111",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"bbb", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"333", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"111", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"444", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ddd", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"ddd",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"222", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"777", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"aaa", x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"222", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"333",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"888", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"eee", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"eee", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"666", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"bbb", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"444", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"444", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"777",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd",
    -- x"000", x"000", x"000", x"000", x"eee", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"444", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"bbb", x"333", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"555",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"444", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"ccc",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"aaa", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"333", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"444", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"222", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"666", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"ccc", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"444", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"777", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ccc", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"777", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"222",
    -- x"000", x"000", x"000", x"111", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"333", x"222", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"888", x"eee", x"fff", x"fff", x"fff",
    -- x"666", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"777",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"444", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"777", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"777", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"ddd", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"eee", x"333", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"eee", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"777", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"888", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"555", x"000",
    -- x"000", x"000", x"000", x"666", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"444", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"333", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"eee", x"222", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"888",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"bbb", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"111", x"666", x"888", x"888",
    -- x"888", x"999", x"bbb", x"ddd", x"fff", x"fff", x"fff", x"eee",
    -- x"ccc", x"777", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"222", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"222", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"999", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"555", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ddd", x"111", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"555", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"444", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"444", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"111", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"666", x"000", x"000",
    -- x"000", x"000", x"000", x"999", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"eee", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"666", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"999", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"aaa",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"666", x"000", x"000", x"000", x"000", x"000", x"000", x"111",
    -- x"555", x"888", x"aaa", x"ddd", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ccc", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"666", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"666", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"555", x"ccc", x"fff", x"fff",
    -- x"ddd", x"444", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"888", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"888", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"eee", x"444", x"000", x"000", x"000",
    -- x"000", x"000", x"444", x"ddd", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"999",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"bbb",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"333", x"000", x"000", x"000", x"666", x"aaa", x"eee", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"777", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"999", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ccc", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"444", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"666", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ddd", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"999",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"888", x"eee", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"666",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"999", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"666",
    -- x"777", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"555", x"222",
    -- x"555", x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"888", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"ddd", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"666", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"333", x"888",
    -- x"222", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"bbb", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"666", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"ccc",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"888", x"555", x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"ccc", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"ddd", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"888", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"999", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"444", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"333", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"666", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"111", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"777",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"555", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"666",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"777", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"111",
    -- x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"888", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"777", x"fff", x"fff",
    -- x"eee", x"222", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"111", x"ccc", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"999", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"eee", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"222", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"555", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"666", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"666", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"444", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"eee", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"444", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"111", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"555", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"777",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"111",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"888", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"000",
    -- x"000", x"333", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"888", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"444", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"999", x"fff", x"fff", x"fff",
    -- x"fff", x"aaa", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"222", x"ddd", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"bbb", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"222", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"888", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"888", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"111", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"222", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ccc", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"222", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"666", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"eee", x"333", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"111", x"aaa", x"eee", x"fff", x"fff",
    -- x"ddd", x"222", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"222", x"999",
    -- x"ddd", x"fff", x"ddd", x"111", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"555", x"bbb",
    -- x"eee", x"fff", x"fff", x"eee", x"888", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"999", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"999", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000",
    -- x"000", x"000", x"999", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"888", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"777", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"888", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"333", x"eee", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"888", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"888", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"222", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"555",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"ddd", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"eee", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ddd", x"111", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"444", x"eee", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"444", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"333", x"aaa", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"666", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"111", x"bbb", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000",
    -- x"000", x"000", x"111", x"eee", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"888",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"333", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"222", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"222", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"555", x"eee", x"fff", x"fff", x"fff", x"fff", x"ddd",
    -- x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"333", x"eee", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"666", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"444", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"888", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"888", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"333", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"bbb",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ccc", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"222", x"eee", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ccc", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"444", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"000", x"000", x"111", x"777", x"bbb", x"ccc", x"bbb",
    -- x"888", x"333", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"222", x"eee", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"666", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"222", x"ddd", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"111", x"ccc", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"444", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"777", x"000",
    -- x"000", x"000", x"000", x"666", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"666", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"eee", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"888", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"777", x"000", x"000", x"000", x"000", x"000",
    -- x"555", x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"000",
    -- x"000", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"888", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"666", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"555", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"666", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"444", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"111",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"999", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"999", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"bbb", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"333", x"ddd", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"333", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"777", x"666", x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"bbb", x"222", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"ccc", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"222", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"111", x"ddd", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"333", x"ddd", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ddd", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"444", x"000",
    -- x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ccc", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"bbb", x"000", x"000", x"000", x"000", x"666",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000",
    -- x"333", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"333", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"888", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"eee", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"888", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"444", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"777", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"555",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"666", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"777", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"aaa", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"111", x"ccc", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"333",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"222", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"888", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"222", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"222", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"666", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"222", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"eee", x"000", x"000", x"000", x"555", x"fff",
    -- x"fff", x"fff", x"fff", x"ccc", x"555", x"000", x"000", x"000",
    -- x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ddd", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"444", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee",
    -- x"ddd", x"bbb", x"aaa", x"999", x"999", x"888", x"666", x"222",
    -- x"000", x"000", x"111", x"555", x"999", x"bbb", x"eee", x"fff",
    -- x"fff", x"fff", x"555", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"777", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"777",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ccc", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"888",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"333", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"eee", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"222", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"666", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"999", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"bbb", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"555", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"444", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"888", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"111", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"eee", x"aaa", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"222", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"111", x"ccc", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"777", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"666", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"888", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"777", x"222", x"bbb", x"fff", x"fff",
    -- x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"000", x"111",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"333", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ccc", x"444", x"111", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"222",
    -- x"555", x"777", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"222", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"aaa", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ddd", x"111", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"aaa",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"bbb", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"999", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"aaa",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"555", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"777", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"333", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"111", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"888", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"111",
    -- x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"444", x"888", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"111", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"aaa",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"444", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"888", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"555", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"999", x"000", x"000", x"000", x"000", x"000", x"999",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"888", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"777", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd",
    -- x"444", x"444", x"555", x"222", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ddd", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"333", x"ddd", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"222", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"bbb",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"ccc", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"555", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"444", x"eee", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"777", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"333",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"888", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ccc", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"777",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"111", x"ccc",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ddd", x"333", x"000", x"aaa", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"444", x"aaa", x"eee", x"fff", x"fff", x"eee", x"bbb", x"555",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"111", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"888", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"999", x"000", x"000", x"000", x"000", x"000", x"222", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"ddd", x"fff", x"fff", x"bbb", x"999", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"555",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"777", x"eee", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"ddd",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"888", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ccc", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"222", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"555", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee",
    -- x"333", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"888", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"555",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"888", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"555", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"111", x"ccc", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc",
    -- x"111", x"000", x"000", x"eee", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"999", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"aaa", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"444", x"ddd", x"fff", x"fff", x"ddd",
    -- x"777", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"222", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"888",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"bbb", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"111",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"555", x"555", x"000", x"000", x"222", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"444", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"222", x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"444", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"888",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"777", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"555", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"333", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"555", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"222", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"444", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"222",
    -- x"888", x"999", x"888", x"444", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"444", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"555", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"111",
    -- x"888", x"ddd", x"fff", x"fff", x"eee", x"999", x"111", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"222", x"ccc", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"000",
    -- x"000", x"000", x"666", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"555", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"555", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"333", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"222", x"eee", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"999", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"777", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"666", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"333", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"555", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"333",
    -- x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"666",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"333", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"888", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"222", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"111", x"ddd", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"eee", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"666", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"222", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"999", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"222",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"333", x"ddd", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"333", x"000",
    -- x"000", x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"eee", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"ddd", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"222", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"444", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"444", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"111", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"555", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"888", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"777", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"666", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"333", x"bbb", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"222", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"333",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"444", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"888",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"eee", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"111", x"ddd", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"222", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"333", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"ccc", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"222", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"aaa", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"555", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"111", x"ddd", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ccc", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"444", x"ddd", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"333", x"eee", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000",
    -- x"000", x"666", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"eee", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"eee", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"777", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"666", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"eee", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"555", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"888", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"333", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"555", x"000", x"000",
    -- x"000", x"000", x"000", x"333", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ddd", x"555", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"444", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"666",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"666", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"222", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"999", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"444",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999",
    -- x"000", x"000", x"000", x"222", x"999", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"222", x"000",
    -- x"000", x"000", x"000", x"000", x"888", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"666", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ddd", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"444", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"666", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"111", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ccc", x"000", x"000", x"000",
    -- x"000", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"111", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"111", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"eee", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000",
    -- x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"777", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"666", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"444", x"000", x"000",
    -- x"000", x"444", x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd",
    -- x"777", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"666", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"ddd",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"111",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"555", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"444", x"111", x"ccc",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"aaa", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"555", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"555", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"000", x"000",
    -- x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"555", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"999", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"333", x"000", x"000", x"000",
    -- x"000", x"000", x"888", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"bbb", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"eee", x"222", x"000", x"000", x"000",
    -- x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"333", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"888",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"999", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"000", x"000",
    -- x"000", x"000", x"444", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"777", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"555", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"999", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"777", x"222", x"777",
    -- x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"666", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"777", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"999", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"777", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000", x"666",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"888", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"888", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"222", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"555", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"333", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"777", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"000", x"000",
    -- x"000", x"000", x"222", x"eee", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"ddd", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"666", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"777", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000",
    -- x"000", x"666", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"111", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"444", x"000", x"000", x"000", x"333",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"eee", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"999", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"555", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"999", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"888", x"000",
    -- x"000", x"222", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"888", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"666", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"666", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"eee", x"aaa", x"333", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"888", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"222", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"666", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"000", x"aaa",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"666", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"bbb",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"666", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"111", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000",
    -- x"000", x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"999", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"666", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000", x"000",
    -- x"333", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"666", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"999",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"666", x"000", x"000", x"000", x"000", x"ddd",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"666", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"999", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"888", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"111",
    -- x"222", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"888", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"888", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"666", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"777", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"999", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"888", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"eee", x"222", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"777", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ddd", x"111", x"000", x"000", x"000", x"000", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"444", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"222",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"888", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"eee", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000",
    -- x"000", x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"666",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"777", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"444",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc",
    -- x"666", x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"444", x"000", x"000", x"000", x"444",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"bbb", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"111", x"888", x"eee", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"888", x"000", x"000", x"000", x"000", x"999", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"333", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"444", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"444",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"777",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"444",
    -- x"ddd", x"fff", x"fff", x"fff", x"fff", x"ddd", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"aaa", x"333",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"bbb", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"555", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"444", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"666", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"888", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"eee", x"222", x"000", x"000", x"000", x"000", x"222", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"777", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"bbb", x"555", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"666", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"111", x"000", x"000",
    -- x"777", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"222",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"333", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"444", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000",
    -- x"000", x"777", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"eee", x"000", x"000", x"000", x"333", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"777", x"eee", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"bbb", x"000", x"000", x"000", x"000", x"555", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"222", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"111", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"777",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"666",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"aaa", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ccc", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"888", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"ccc", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"888", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ccc", x"777", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"ccc", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"333", x"ddd", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee",
    -- x"333", x"000", x"000", x"000", x"000", x"000", x"000", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"000",
    -- x"444", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"555", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"444",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"444", x"eee", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000", x"000",
    -- x"000", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"ddd", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"555", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"888", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee",
    -- x"111", x"000", x"000", x"000", x"222", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"eee", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"999",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"444",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"999", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"eee", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"333", x"ccc", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"333", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"555", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"aaa", x"333", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"ddd", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"111", x"ddd", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"999",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"444",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"777", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"666",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"bbb", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"333", x"000", x"333", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"888", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000", x"000",
    -- x"000", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"444", x"000", x"000", x"999", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"bbb", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"777", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"777",
    -- x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ccc", x"bbb", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"444", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"111", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ccc", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"bbb",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"888", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"222", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ccc", x"000", x"000", x"000", x"000", x"999",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"111",
    -- x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"999",
    -- x"111", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"ddd", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"333", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"999", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"444", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"ddd",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"111", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"aaa", x"000", x"000", x"222", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"444", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"444", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"999", x"000", x"333", x"eee", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"444",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"222", x"000",
    -- x"000", x"000", x"000", x"333", x"eee", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"000",
    -- x"666", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ccc", x"000", x"000", x"999", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ccc", x"444", x"111", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"222", x"000", x"000", x"000", x"000",
    -- x"555", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"000",
    -- x"000", x"000", x"000", x"aaa", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"bbb", x"000", x"333", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"666", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"ccc",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"555", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"333", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ddd", x"111", x"000", x"000", x"000", x"000", x"111",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ccc", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"111", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"444", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"999",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"bbb", x"333", x"111", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"eee", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"666", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"eee", x"333", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"777",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"222", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"bbb", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"eee", x"000", x"000", x"ccc", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"eee", x"aaa", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"222", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000",
    -- x"000", x"000", x"000", x"ccc", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"bbb", x"000", x"000", x"000", x"000", x"000",
    -- x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"777", x"000", x"999", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"777", x"000", x"000", x"000", x"555",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000", x"000",
    -- x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"333", x"000",
    -- x"000", x"000", x"777", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"666", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"999", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"ddd",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"888", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ddd", x"111", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"eee", x"111", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"555",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"888", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"555", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"888", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"222", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"eee", x"333", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"111", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"333",
    -- x"000", x"000", x"000", x"000", x"000", x"777", x"aaa", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"ccc", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"eee", x"777", x"ddd", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"999", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"555", x"333", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"eee", x"333", x"333", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"ddd", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd",
    -- x"bbb", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"aaa", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"000", x"777", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"555", x"000", x"000", x"000", x"000", x"000",
    -- x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"777", x"999", x"eee",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000", x"000",
    -- x"000", x"555", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee",
    -- x"111", x"000", x"000", x"000", x"888", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"111",
    -- x"000", x"000", x"000", x"000", x"000", x"888", x"aaa", x"000",
    -- x"000", x"000", x"000", x"ccc", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"666", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"555", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999",
    -- x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"555", x"ddd",
    -- x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd",
    -- x"111", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"222", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ccc", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"777", x"ddd", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ddd", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"555", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"666", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"222", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"999",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"222", x"999", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ddd", x"222", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"555", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"000",
    -- x"000", x"000", x"000", x"000", x"888", x"fff", x"fff", x"222",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"777", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ccc", x"111", x"000", x"bbb", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"444",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"777", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"333", x"000", x"000", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"888", x"aaa", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"777", x"000", x"000", x"000", x"000", x"000", x"000", x"333",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ddd", x"444", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ddd", x"333", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"eee", x"111", x"000", x"000",
    -- x"444", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"666",
    -- x"000", x"000", x"000", x"000", x"333", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc",
    -- x"222", x"000", x"000", x"222", x"bbb", x"fff", x"fff", x"111",
    -- x"000", x"000", x"000", x"ddd", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"444", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"111", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"555", x"fff", x"fff", x"fff", x"fff", x"ddd", x"333", x"000",
    -- x"000", x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"333", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"777", x"fff", x"fff",
    -- x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"111",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"444", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"222",
    -- x"bbb", x"fff", x"fff", x"777", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"999", x"eee", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"444", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"444", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"999", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"111",
    -- x"777", x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ddd", x"111", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"888", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000",
    -- x"000", x"000", x"111", x"bbb", x"fff", x"fff", x"fff", x"999",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"777",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"999", x"000", x"000", x"000", x"eee", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"444", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"eee", x"333", x"000", x"000", x"000", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000",
    -- x"000", x"000", x"000", x"000", x"888", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"aaa", x"000", x"111", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"666",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"999",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb",
    -- x"111", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"222", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"666", x"000", x"000", x"333",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ccc", x"ddd", x"fff", x"fff", x"fff", x"fff", x"999",
    -- x"000", x"000", x"000", x"ddd", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"333", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"ddd", x"fff", x"fff", x"ccc", x"111", x"000", x"000",
    -- x"000", x"222", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"999", x"fff", x"fff", x"fff",
    -- x"ddd", x"ddd", x"fff", x"fff", x"fff", x"bbb", x"111", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"777", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"222", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"666", x"eee",
    -- x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ddd", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"111", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"333", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"666", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"999", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"111", x"000",
    -- x"000", x"000", x"000", x"444", x"888", x"aaa", x"ddd", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ddd", x"111", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"aaa", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"888", x"000",
    -- x"000", x"333", x"ddd", x"fff", x"fff", x"fff", x"fff", x"eee",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"888", x"888", x"111", x"000", x"ddd",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"777", x"000", x"000", x"000", x"333", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"111", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"888", x"000", x"000", x"000", x"000", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"000",
    -- x"000", x"000", x"000", x"666", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ccc", x"000", x"000", x"000", x"bbb", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"eee", x"fff", x"666", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"ccc",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"777", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"555", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"333", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"555", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee",
    -- x"000", x"000", x"000", x"eee", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"eee", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"666", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"999", x"fff", x"ccc", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"888", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"000", x"000",
    -- x"000", x"000", x"444", x"ccc", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"bbb", x"fff", x"fff", x"666", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"444",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ddd", x"333", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"333", x"bbb", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"555", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"eee", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"eee", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"777", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"eee", x"222", x"000", x"555",
    -- x"999", x"ccc", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"222", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"ccc", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"666", x"000",
    -- x"777", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"777", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"111", x"888", x"eee", x"fff", x"fff", x"999", x"000", x"ccc",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"000", x"000", x"000", x"000", x"777", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"111",
    -- x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"222", x"000", x"000", x"000", x"000", x"ddd", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"000",
    -- x"000", x"000", x"777", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ddd", x"111", x"000", x"000", x"000", x"666", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"222", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"444", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"ccc", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"777", x"000", x"444", x"eee", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"555", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"666", x"000", x"000", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ccc", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"888", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"222", x"ccc", x"111", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"ccc", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"aaa",
    -- x"bbb", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ccc", x"ddd", x"333", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"444", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"666",
    -- x"888", x"aaa", x"bbb", x"ddd", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ccc", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"ddd", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"888", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"444", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"eee", x"888", x"bbb", x"eee", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"eee", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"666", x"bbb",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee",
    -- x"444", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"222", x"999",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"888", x"666", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"999",
    -- x"222", x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"333", x"ddd",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb",
    -- x"111", x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"111",
    -- x"555", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee",
    -- x"333", x"000", x"000", x"000", x"000", x"000", x"ddd", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"999", x"111", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"777", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"999", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"111", x"888", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"ddd", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee",
    -- x"333", x"000", x"000", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"bbb", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"aaa", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"222", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"333", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"888", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"444", x"eee", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"ddd", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"eee", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"888", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ccc", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"222", x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"666", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"111", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc", x"222",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"222", x"aaa", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"777", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"ddd",
    -- x"bbb", x"aaa", x"999", x"777", x"444", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"555",
    -- x"000", x"000", x"000", x"000", x"111", x"999", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"555",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"555", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"bbb", x"333", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"bbb", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ccc", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"666", x"000", x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"111", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"555", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"333",
    -- x"000", x"000", x"222", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"999", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"ccc", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"666", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"eee", x"999", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"555", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"111", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"eee", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"555", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"444", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"777", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ccc", x"777", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"555", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"333", x"aaa", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"eee", x"777", x"888", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"aaa", x"aaa", x"ccc", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"eee", x"666", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"888", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"888", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"777",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"555", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"111", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ddd", x"111", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"333", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"333",
    -- x"000", x"000", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"eee", x"222", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"aaa",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"444", x"000",
    -- x"000", x"000", x"555", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"777", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"eee", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"888", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"444",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ddd", x"333", x"000", x"777", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ddd", x"444", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"444", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"999", x"fff", x"fff",
    -- x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"444", x"ccc",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"888", x"333", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"888", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"444", x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"bbb", x"222", x"bbb", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"bbb", x"999", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ccc", x"222", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"555", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"333", x"bbb", x"eee", x"fff", x"fff", x"fff", x"bbb", x"555",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"777", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"333", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"666", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"111", x"000",
    -- x"000", x"555", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"444", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"666", x"000", x"000",
    -- x"000", x"000", x"888", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"555", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"222", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"555", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"111", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"111", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"888", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ddd", x"111", x"000", x"000", x"000", x"777", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"999", x"111", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"666", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"999", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff",
    -- x"fff", x"eee", x"222", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"999", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"ddd", x"ddd", x"ccc", x"aaa", x"666", x"111",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"888", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"444", x"bbb",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"777", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"555", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"bbb", x"000", x"000", x"999", x"eee", x"fff",
    -- x"fff", x"ccc", x"666", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"111", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"222", x"444", x"111", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"eee", x"444", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"444", x"bbb",
    -- x"eee", x"fff", x"fff", x"ccc", x"666", x"000", x"000", x"000",
    -- x"000", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"555", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"777", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"666", x"000", x"000", x"000",
    -- x"000", x"000", x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"444", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"666", x"fff", x"fff",
    -- x"fff", x"fff", x"ddd", x"555", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"999", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd",
    -- x"111", x"000", x"000", x"000", x"000", x"000", x"777", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"999", x"222",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"555", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"444", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"ccc", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"eee", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ddd", x"fff", x"fff",
    -- x"fff", x"666", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"444", x"999", x"ddd", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"eee", x"999", x"888", x"666", x"444",
    -- x"111", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"777", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"333", x"bbb", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"666", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"ccc", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"aaa", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"ddd", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ccc", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"111", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"555", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"666", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"666", x"aaa", x"ccc", x"ddd", x"eee",
    -- x"ddd", x"ccc", x"999", x"222", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"111", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff",
    -- x"fff", x"ccc", x"111", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"111", x"eee", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ddd", x"444", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"222",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"777",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"eee", x"888", x"111", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"333", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"111", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"666", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"999", x"fff", x"fff",
    -- x"bbb", x"000", x"000", x"000", x"000", x"000", x"222", x"888",
    -- x"bbb", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ccc", x"222", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"666", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ddd", x"444", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"444", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee",
    -- x"666", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"999", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ddd", x"111", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"555",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"555", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"888",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"999", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"eee", x"fff", x"fff",
    -- x"ddd", x"111", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"666", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"999", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"777",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"333", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"666", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"888", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"222", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"333", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"333", x"fff", x"bbb",
    -- x"000", x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"999", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"333", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"999", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"777", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb",
    -- x"111", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"666",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"999", x"111",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"111", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ccc", x"222", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"666", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"888", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"666", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"bbb", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"444", x"fff", x"fff", x"eee",
    -- x"333", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"333",
    -- x"999", x"ccc", x"eee", x"fff", x"fff", x"fff", x"eee", x"aaa",
    -- x"222", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"111", x"fff",
    -- x"fff", x"fff", x"fff", x"eee", x"999", x"222", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"555", x"bbb", x"eee", x"fff", x"fff", x"fff", x"ccc",
    -- x"888", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"555", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee",
    -- x"555", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ccc",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"444", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"888", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"444", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"888", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"555",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"aaa", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"777", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"888", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ddd", x"222", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"222", x"fff", x"ddd", x"333",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"111", x"eee",
    -- x"fff", x"ccc", x"777", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"eee", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"666", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"aaa", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"111",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"111",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ddd", x"333", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"888", x"ccc", x"fff", x"fff", x"eee", x"ccc",
    -- x"bbb", x"888", x"333", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"333", x"bbb", x"eee", x"fff", x"fff", x"eee", x"aaa", x"333",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"999", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"777", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"555", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"aaa", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"999", x"fff", x"ddd", x"aaa", x"777", x"333",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"111", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"eee", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"555", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"777", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ccc", x"444", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"333", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"888", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"eee", x"888", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"666", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"444", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"333", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"444", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ddd", x"666", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"ccc", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"444", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"aaa", x"222", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"111", x"ccc", x"fff", x"fff",
    -- x"eee", x"ccc", x"444", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"666", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"eee", x"555", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"111", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"999", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"222", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"666", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"666", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa",
    -- x"333", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"555", x"ccc", x"eee", x"fff", x"fff", x"ddd",
    -- x"888", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"eee", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"bbb", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"aaa", x"111",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"111", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"222", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"888", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"eee", x"999", x"222", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ddd", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"333", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"333", x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ddd", x"999", x"333", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"aaa", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"111", x"999", x"ddd", x"fff",
    -- x"fff", x"ddd", x"aaa", x"555", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ccc", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ccc", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"444", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"666", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"333", x"ddd", x"fff", x"fff", x"eee", x"ccc", x"aaa",
    -- x"888", x"555", x"111", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"555", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"222", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"111",
    -- x"222", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"aaa", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"777", x"eee", x"fff", x"ccc",
    -- x"555", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"333", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"111",
    -- x"eee", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"aaa", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"333", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"333", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"aaa",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"222", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"555", x"ddd",
    -- x"fff", x"fff", x"aaa", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"777", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"444", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"888", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"ddd", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"222", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"666", x"999",
    -- x"999", x"999", x"888", x"888", x"777", x"777", x"666", x"666",
    -- x"666", x"555", x"555", x"555", x"555", x"555", x"555", x"444",
    -- x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444",
    -- x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444",
    -- x"444", x"444", x"444", x"444", x"444", x"555", x"555", x"666",
    -- x"666", x"777", x"888", x"999", x"999", x"999", x"555", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"777",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"ddd", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"bbb", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"777", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"444",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"999", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"ddd", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"eee", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"444", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"666", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"999", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"222", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"888", x"ddd", x"ccc", x"ccc", x"bbb", x"bbb",
    -- x"aaa", x"999", x"999", x"999", x"999", x"888", x"888", x"888",
    -- x"888", x"999", x"999", x"999", x"999", x"aaa", x"aaa", x"aaa",
    -- x"bbb", x"bbb", x"bbb", x"ccc", x"ccc", x"ccc", x"ddd", x"ddd",
    -- x"ddd", x"eee", x"eee", x"eee", x"eee", x"eee", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"111",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"555", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"bbb", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"ccc", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"444", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"222", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"ccc", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"999", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"555", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"ddd", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"ccc", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"111",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"fff", x"555", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"666",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"ddd", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"999",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"fff", x"666", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"ccc",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"ddd", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"eee",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"fff", x"555", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"222", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"ccc", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"444", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff",
    -- x"333", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"666", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"999",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"888", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"ddd", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"777", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"fff", x"444", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"444", x"fff",
    -- x"fff", x"fff", x"fff", x"fff", x"fff", x"666", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"aaa",
    -- x"eee", x"fff", x"fff", x"ddd", x"555", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000",
    -- x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"
-- );
 
 
end package;